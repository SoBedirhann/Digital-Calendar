`timescale 1ns / 1ps

module char_rom(
    input wire [3:0] char_code, // Gösterilecek karakterin kodu (0-9, A-F)
    input wire [4:0] row,       // Karakterin sat?r indeksi (0-7)
    output reg [31:0] pixel_row  // Karakterin o sat?rdaki piksel verisi
);

    // Karakter ROM'u (her karakter 8x8 bit)
    always @* begin
        case (char_code)
            4'h0: begin
            // " 0 "
                case (row)
                    5'd0:  pixel_row = 32'b00000000011111111111111100000000;
                    5'd1:  pixel_row = 32'b00000001111111111111111110000000;
                    5'd2:  pixel_row = 32'b00000011111000000000111111000000;
                    5'd3:  pixel_row = 32'b00000111110000000000011111100000;
                    5'd4:  pixel_row = 32'b00001111100000000000001111110000;
                    5'd5:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd6:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd7:  pixel_row = 32'b00111110000000000000000011111100;
                    5'd8:  pixel_row = 32'b00111110000000000000000011111100;
                    5'd9:  pixel_row = 32'b00111110000000000000000011111100;
                    5'd10: pixel_row = 32'b01111100000000000000000001111110;
                    5'd11: pixel_row = 32'b01111100000000000000000001111110;
                    5'd12: pixel_row = 32'b01111100000000000000000001111110;
                    5'd13: pixel_row = 32'b01111100000000000000000001111110;
                    5'd14: pixel_row = 32'b01111100000000000000000001111110;
                    5'd15: pixel_row = 32'b01111100000000000000000001111110;
                    5'd16: pixel_row = 32'b01111100000000000000000001111110;
                    5'd17: pixel_row = 32'b01111100000000000000000001111110;
                    5'd18: pixel_row = 32'b01111100000000000000000001111110;
                    5'd19: pixel_row = 32'b01111100000000000000000001111110;
                    5'd20: pixel_row = 32'b01111100000000000000000001111110;
                    5'd21: pixel_row = 32'b01111100000000000000000001111110;
                    5'd22: pixel_row = 32'b00111110000000000000000011111100;
                    5'd23: pixel_row = 32'b00111110000000000000000011111100;
                    5'd24: pixel_row = 32'b00111110000000000000000011111100;
                    5'd25: pixel_row = 32'b00011111000000000000000111111000;
                    5'd26: pixel_row = 32'b00011111000000000000000111111000;
                    5'd27: pixel_row = 32'b00001111100000000000001111110000;
                    5'd28: pixel_row = 32'b00000111110000000000011111100000;
                    5'd29: pixel_row = 32'b00000011111000000000111111000000;
                    5'd30: pixel_row = 32'b00000001111111111111111110000000;
                    5'd31: pixel_row = 32'b00000000011111111111111100000000;
                endcase
            end
            4'h1: begin
            // " 1 "
                case (row)
                    5'd0:  pixel_row = 32'b00000000000011111100000000000000;
                    5'd1:  pixel_row = 32'b00000000000111111100000000000000;
                    5'd2:  pixel_row = 32'b00000000001111111100000000000000;
                    5'd3:  pixel_row = 32'b00000000011111111100000000000000;
                    5'd4:  pixel_row = 32'b00000000111101111100000000000000;
                    5'd5:  pixel_row = 32'b00000000111001111100000000000000;
                    5'd6:  pixel_row = 32'b00000001110001111100000000000000;
                    5'd7:  pixel_row = 32'b00000001100001111100000000000000;
                    5'd8:  pixel_row = 32'b00000011000001111100000000000000;
                    5'd9:  pixel_row = 32'b00000011000001111100000000000000;
                    5'd10: pixel_row = 32'b00000000000001111100000000000000;
                    5'd11: pixel_row = 32'b00000000000001111100000000000000;
                    5'd12: pixel_row = 32'b00000000000001111100000000000000;
                    5'd13: pixel_row = 32'b00000000000001111100000000000000;
                    5'd14: pixel_row = 32'b00000000000001111100000000000000;
                    5'd15: pixel_row = 32'b00000000000001111100000000000000;
                    5'd16: pixel_row = 32'b00000000000001111100000000000000;
                    5'd17: pixel_row = 32'b00000000000001111100000000000000;
                    5'd18: pixel_row = 32'b00000000000001111100000000000000;
                    5'd19: pixel_row = 32'b00000000000001111100000000000000;
                    5'd20: pixel_row = 32'b00000000000001111100000000000000;
                    5'd21: pixel_row = 32'b00000000000001111100000000000000;
                    5'd22: pixel_row = 32'b00000000000001111100000000000000;
                    5'd23: pixel_row = 32'b00000000000001111100000000000000;
                    5'd24: pixel_row = 32'b00000000000001111100000000000000;
                    5'd25: pixel_row = 32'b00000000000001111100000000000000;
                    5'd26: pixel_row = 32'b00000000000001111100000000000000;
                    5'd27: pixel_row = 32'b00000000000001111100000000000000;
                    5'd28: pixel_row = 32'b00000000000001111100000000000000;
                    5'd29: pixel_row = 32'b11111111111111111111111111111100;
                    5'd30: pixel_row = 32'b11111111111111111111111111111100;
                    5'd31: pixel_row = 32'b11111111111111111111111111111100;
                endcase
            end
            4'h2: begin
            // " 2 "
                case (row)
                    5'd0:  pixel_row = 32'b00000000011111111111111100000000;
                    5'd1:  pixel_row = 32'b00000001111111111111111110000000;
                    5'd2:  pixel_row = 32'b00000011111100000000111111000000;
                    5'd3:  pixel_row = 32'b00000111110000000000011111100000;
                    5'd4:  pixel_row = 32'b00001111100000000000001111110000;
                    5'd5:  pixel_row = 32'b00001111100000000000001111110000;
                    5'd6:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd7:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd8:  pixel_row = 32'b00000000000000000000000111111000;
                    5'd9:  pixel_row = 32'b00000000000000000000000111111000;
                    5'd10: pixel_row = 32'b00000000000000000000000111110000;
                    5'd11: pixel_row = 32'b00000000000000000000001111110000;
                    5'd12: pixel_row = 32'b00000000000000000000011111100000;
                    5'd13: pixel_row = 32'b00000000000000000000111111000000;
                    5'd14: pixel_row = 32'b00000000000000000001111110000000;
                    5'd15: pixel_row = 32'b00000000000000000011111100000000;
                    5'd16: pixel_row = 32'b00000000000000000111111000000000;
                    5'd17: pixel_row = 32'b00000000000000001111110000000000;
                    5'd18: pixel_row = 32'b00000000000000011111100000000000;
                    5'd19: pixel_row = 32'b00000000000000111111000000000000;
                    5'd20: pixel_row = 32'b00000000000001111110000000000000;
                    5'd21: pixel_row = 32'b00000000000011111100000000000000;
                    5'd22: pixel_row = 32'b00000000000111111000000000000000;
                    5'd23: pixel_row = 32'b00000000001111110000000000000000;
                    5'd24: pixel_row = 32'b00000000011111100000000000000000;
                    5'd25: pixel_row = 32'b00000000111111000000000000000000;
                    5'd26: pixel_row = 32'b00000001111110000000000000000000;
                    5'd27: pixel_row = 32'b00000011111100000000000000000000;
                    5'd28: pixel_row = 32'b00000111111111111111111111111100;
                    5'd29: pixel_row = 32'b00001111111111111111111111111100;
                    5'd30: pixel_row = 32'b00011111111111111111111111111100;
                    5'd31: pixel_row = 32'b11111111111111111111111111111100;
                endcase
            end
            4'h3: begin
            // " 3 "
                case (row)
                    5'd0:  pixel_row = 32'b00000000011111111111111100000000;
                    5'd1:  pixel_row = 32'b00000001111111111111111110000000;
                    5'd2:  pixel_row = 32'b00000011111100000000111111000000;
                    5'd3:  pixel_row = 32'b00000111110000000000011111100000;
                    5'd4:  pixel_row = 32'b00001111100000000000001111110000;
                    5'd5:  pixel_row = 32'b00001111100000000000001111110000;
                    5'd6:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd7:  pixel_row = 32'b00011111000000000000000111111000;
                    5'd8:  pixel_row = 32'b00000000000000000000000111111000;
                    5'd9:  pixel_row = 32'b00000000000000000000000111111000;
                    5'd10: pixel_row = 32'b00000000000000000000000111110000;
                    5'd11: pixel_row = 32'b00000000000000000000011111100000;
                    5'd12: pixel_row = 32'b00000000000000001111111110000000;
                    5'd13: pixel_row = 32'b00000000000000011111111100000000;
                    5'd14: pixel_row = 32'b00000000000000000000011111000000;
                    5'd15: pixel_row = 32'b00000000000000000000001111110000;
                    5'd16: pixel_row = 32'b00000000000000000000000111111000;
                    5'd17: pixel_row = 32'b00000000000000000000000111111000;
                    5'd18: pixel_row = 32'b00000000000000000000000111111000;
                    5'd19: pixel_row = 32'b00000000000000000000000111111000;
                    5'd20: pixel_row = 32'b00000000000000000000000111111000;
                    5'd21: pixel_row = 32'b00000000000000000000000111111000;
                    5'd22: pixel_row = 32'b00011111000000000000000111111000;
                    5'd23: pixel_row = 32'b00011111000000000000000111111000;
                    5'd24: pixel_row = 32'b00001111100000000000001111110000;
                    5'd25: pixel_row = 32'b00001111100000000000001111110000;
                    5'd26: pixel_row = 32'b00000111110000000000011111100000;
                    5'd27: pixel_row = 32'b00000011111100000000111111000000;
                    5'd28: pixel_row = 32'b00000001111111111111111110000000;
                    5'd29: pixel_row = 32'b00000000011111111111111100000000;
                    5'd30: pixel_row = 32'b00000000000000000000000000000000;
                    5'd31: pixel_row = 32'b00000000000000000000000000000000;
                endcase
            end
            4'hA: begin 
            // ':' karakteri için
                case (row)
                    5'd0:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd1:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd2:  pixel_row = 32'b00000000000000001111100000000000;
                    5'd3:  pixel_row = 32'b00000000000000011111110000000000;
                    5'd4:  pixel_row = 32'b00000000000000111111111000000000;
                    5'd5:  pixel_row = 32'b00000000000000111111111000000000;
                    5'd6:  pixel_row = 32'b00000000000000011111110000000000;
                    5'd7:  pixel_row = 32'b00000000000000001111100000000000;
                    5'd8:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd9:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd10: pixel_row = 32'b00000000000000000000000000000000;
                    5'd11: pixel_row = 32'b00000000000000000000000000000000;
                    5'd12: pixel_row = 32'b00000000000000000000000000000000;
                    5'd13: pixel_row = 32'b00000000000000000000000000000000;
                    5'd14: pixel_row = 32'b00000000000000000000000000000000;
                    5'd15: pixel_row = 32'b00000000000000000000000000000000;
                    5'd16: pixel_row = 32'b00000000000000000000000000000000;
                    5'd17: pixel_row = 32'b00000000000000000000000000000000;
                    5'd18: pixel_row = 32'b00000000000000001111100000000000;
                    5'd19: pixel_row = 32'b00000000000000011111110000000000;
                    5'd20: pixel_row = 32'b00000000000000111111111000000000;
                    5'd21: pixel_row = 32'b00000000000000111111111000000000;
                    5'd22: pixel_row = 32'b00000000000000011111110000000000;
                    5'd23: pixel_row = 32'b00000000000000001111100000000000;
                    5'd24: pixel_row = 32'b00000000000000000000000000000000;
                    5'd25: pixel_row = 32'b00000000000000000000000000000000;
                    5'd26: pixel_row = 32'b00000000000000000000000000000000;
                    5'd27: pixel_row = 32'b00000000000000000000000000000000;
                    5'd28: pixel_row = 32'b00000000000000000000000000000000;
                    5'd29: pixel_row = 32'b00000000000000000000000000000000;
                    5'd30: pixel_row = 32'b00000000000000000000000000000000;
                    5'd31: pixel_row = 32'b00000000000000000000000000000000;
                endcase
            end
            4'hB: begin 
            // '.' karakteri için (Bo?luk)
                case (row)
                    5'd0:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd1:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd2:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd3:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd4:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd5:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd6:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd7:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd8:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd9:  pixel_row = 32'b00000000000000000000000000000000;
                    5'd10: pixel_row = 32'b00000000000000000000000000000000;
                    5'd11: pixel_row = 32'b00000000000000000000000000000000;
                    5'd12: pixel_row = 32'b00000000000000000000000000000000;
                    5'd13: pixel_row = 32'b00000000000000000000000000000000;
                    5'd14: pixel_row = 32'b00000000000000000000000000000000;
                    5'd15: pixel_row = 32'b00000000000000000000000000000000;
                    5'd16: pixel_row = 32'b00000000000000000000000000000000;
                    5'd17: pixel_row = 32'b00000000000000000000000000000000;
                    5'd18: pixel_row = 32'b00000000000000001111100000000000;
                    5'd19: pixel_row = 32'b00000000000000011111110000000000;
                    5'd20: pixel_row = 32'b00000000000000111111111000000000;
                    5'd21: pixel_row = 32'b00000000000000111111111000000000;
                    5'd22: pixel_row = 32'b00000000000000011111110000000000;
                    5'd23: pixel_row = 32'b00000000000000001111100000000000;
                    5'd24: pixel_row = 32'b00000000000000000000000000000000;
                    5'd25: pixel_row = 32'b00000000000000000000000000000000;
                    5'd26: pixel_row = 32'b00000000000000000000000000000000;
                    5'd27: pixel_row = 32'b00000000000000000000000000000000;
                    5'd28: pixel_row = 32'b00000000000000000000000000000000;
                    5'd29: pixel_row = 32'b00000000000000000000000000000000;
                    5'd30: pixel_row = 32'b00000000000000000000000000000000;
                    5'd31: pixel_row = 32'b00000000000000000000000000000000;
                endcase
           end
            4'h4: begin // 4 karakteri için
                case (row)
                    5'd0:  pixel_row = 32'b00000000000000000000111100000000;
                    5'd1:  pixel_row = 32'b00000000000000000001111100000000;
                    5'd2:  pixel_row = 32'b00000000000000000011111100000000;
                    5'd3:  pixel_row = 32'b00000000000000000111111100000000;
                    5'd4:  pixel_row = 32'b00000000000000001111111100000000;
                    5'd5:  pixel_row = 32'b00000000000000011111011100000000;
                    5'd6:  pixel_row = 32'b00000000000000111110011100000000;
                    5'd7:  pixel_row = 32'b00000000000001111100011100000000;
                    5'd8:  pixel_row = 32'b00000000000011111000011100000000;
                    5'd9:  pixel_row = 32'b00000000000111110000011100000000;
                    5'd10: pixel_row = 32'b00000000001111100000011100000000;
                    5'd11: pixel_row = 32'b00000000011111000000011100000000;
                    5'd12: pixel_row = 32'b00000000111110000000011100000000;
                    5'd13: pixel_row = 32'b00000001111100000000011100000000;
                    5'd14: pixel_row = 32'b00000011111000000000011100000000;
                    5'd15: pixel_row = 32'b00000111110000000000011100000000;
                    5'd16: pixel_row = 32'b00001111100000000000011100000000;
                    5'd17: pixel_row = 32'b00011111111111111111111111111000;
                    5'd18: pixel_row = 32'b00011111111111111111111111111000;
                    5'd19: pixel_row = 32'b00011111111111111111111111111000;
                    5'd20: pixel_row = 32'b00000000000000000000011100000000;
                    5'd21: pixel_row = 32'b00000000000000000000011100000000;
                    5'd22: pixel_row = 32'b00000000000000000000011100000000;
                    5'd23: pixel_row = 32'b00000000000000000000011100000000;
                    5'd24: pixel_row = 32'b00000000000000000000011100000000;
                    5'd25: pixel_row = 32'b00000000000000000000011100000000;
                    5'd26: pixel_row = 32'b00000000000000000000011100000000;
                    5'd27: pixel_row = 32'b00000000000000000000011100000000;
                    5'd28: pixel_row = 32'b00000000000000000000011100000000;
                    5'd29: pixel_row = 32'b00000000000000000000011100000000;
                    5'd30: pixel_row = 32'b00000000000000000000011100000000;
                    5'd31: pixel_row = 32'b00000000000000000000000000000000;
                endcase
            end
            
            4'h5: begin // 5 karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00000000011111111111111111111000;
        5'd1:  pixel_row = 32'b00000000111111111111111111111000;
        5'd2:  pixel_row = 32'b00000000111111111111111111111000;
        5'd3:  pixel_row = 32'b00000000111111111111111111111000;
        5'd4:  pixel_row = 32'b00000000111100000000000000000000;
        5'd5:  pixel_row = 32'b00000000111100000000000000000000;
        5'd6:  pixel_row = 32'b00000000111100000000000000000000;
        5'd7:  pixel_row = 32'b00000000111100000000000000000000;
        5'd8:  pixel_row = 32'b00000000111100000000000000000000;
        5'd9:  pixel_row = 32'b00000000111100000000000000000000;
        5'd10: pixel_row = 32'b00000000111100000000000000000000;
        5'd11: pixel_row = 32'b00000000111100000000000000000000;
        5'd12: pixel_row = 32'b00000000111100000000000000000000;
        5'd13: pixel_row = 32'b00000000111100000000000000000000;
        5'd14: pixel_row = 32'b00000000111111111111111110000000;
        5'd15: pixel_row = 32'b00000000111111111111111111100000;
        5'd16: pixel_row = 32'b00000000000000000000000111110000;
        5'd17: pixel_row = 32'b00000000000000000000000011111000;
        5'd18: pixel_row = 32'b00000000000000000000000011111000;
        5'd19: pixel_row = 32'b00000000000000000000000001111000;
        5'd20: pixel_row = 32'b00000000000000000000000001111000;
        5'd21: pixel_row = 32'b00000000000000000000000001111000;
        5'd22: pixel_row = 32'b00000000000000000000000001111000;
        5'd23: pixel_row = 32'b00000000000000000000000001111000;
        5'd24: pixel_row = 32'b11110000000000000000000011110000;
        5'd25: pixel_row = 32'b11110000000000000000000011110000;
        5'd26: pixel_row = 32'b01111000000000000000000111100000;
        5'd27: pixel_row = 32'b01111100000000000000011111100000;
        5'd28: pixel_row = 32'b00111111111111111111111111000000;
        5'd29: pixel_row = 32'b00011111111111111111111110000000;
        5'd30: pixel_row = 32'b00000000000000000000000000000000;
        5'd31: pixel_row = 32'b00000000000000000000000000000000;
    endcase
end
            
            4'h6: begin // 6 karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00000000000001111111111110000000;
        5'd1:  pixel_row = 32'b00000000000011111111111111000000;
        5'd2:  pixel_row = 32'b00000000000111111111111111100000;
        5'd3:  pixel_row = 32'b00000000001111100000001111110000;
        5'd4:  pixel_row = 32'b00000000011111000000000011111000;
        5'd5:  pixel_row = 32'b00000000111110000000000011111000;
        5'd6:  pixel_row = 32'b00000001111100000000000011111000;
        5'd7:  pixel_row = 32'b00000001111100000000000011110000;
        5'd8:  pixel_row = 32'b00000011111000000000000000000000;
        5'd9:  pixel_row = 32'b00000111110000000000000000000000;
        5'd10: pixel_row = 32'b00000111100000000000000000000000;
        5'd11: pixel_row = 32'b00001111100000000000000000000000;
        5'd12: pixel_row = 32'b00001111100000000000000000000000;
        5'd13: pixel_row = 32'b00001111000000000000000000000000;
        5'd14: pixel_row = 32'b00011111000000000000000000000000;
        5'd15: pixel_row = 32'b00011111001111111111111000000000;
        5'd16: pixel_row = 32'b00111111111111111111111110000000;
        5'd17: pixel_row = 32'b00111111111111111111111111000000;
        5'd18: pixel_row = 32'b00111111111100000000011111100000;
        5'd19: pixel_row = 32'b00111111110000000000000111100000;
        5'd20: pixel_row = 32'b00111111000000000000000011110000;
        5'd21: pixel_row = 32'b00111110000000000000000011110000;
        5'd22: pixel_row = 32'b00111110000000000000000011110000;
        5'd23: pixel_row = 32'b00111100000000000000000011110000;
        5'd24: pixel_row = 32'b00111100000000000000000011110000;
        5'd25: pixel_row = 32'b00111100000000000000000011110000;
        5'd26: pixel_row = 32'b00111100000000000000000011110000;
        5'd27: pixel_row = 32'b00011110000000000000000111100000;
        5'd28: pixel_row = 32'b00011111000000000000001111100000;
        5'd29: pixel_row = 32'b00001111100000000000011111100000;
        5'd30: pixel_row = 32'b00000111111111111111111111000000;
        5'd31: pixel_row = 32'b00000011111111111111111110000000;
    endcase
end

            4'h7: begin // 7 karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00011111111111111111111111111100;
        5'd1:  pixel_row = 32'b00011111111111111111111111111100;
        5'd2:  pixel_row = 32'b00011111111111111111111111111100;
        5'd3:  pixel_row = 32'b00000000000000000000000111111000;
        5'd4:  pixel_row = 32'b00000000000000000000001111110000;
        5'd5:  pixel_row = 32'b00000000000000000000001111110000;
        5'd6:  pixel_row = 32'b00000000000000000000011111100000;
        5'd7:  pixel_row = 32'b00000000000000000000111111000000;
        5'd8:  pixel_row = 32'b00000000000000000001111110000000;
        5'd9:  pixel_row = 32'b00000000000000000011111100000000;
        5'd10: pixel_row = 32'b00000000000000000011111000000000;
        5'd11: pixel_row = 32'b00000000000000000111110000000000;
        5'd12: pixel_row = 32'b00000000000000001111100000000000;
        5'd13: pixel_row = 32'b00000000000000001111100000000000;
        5'd14: pixel_row = 32'b00000000000000011111000000000000;
        5'd15: pixel_row = 32'b00000000000000111110000000000000;
        5'd16: pixel_row = 32'b00000000000001111100000000000000;
        5'd17: pixel_row = 32'b00000000000001111100000000000000;
        5'd18: pixel_row = 32'b00000000000011111000000000000000;
        5'd19: pixel_row = 32'b00000000000111110000000000000000;
        5'd20: pixel_row = 32'b00000000000111100000000000000000;
        5'd21: pixel_row = 32'b00000000001111100000000000000000;
        5'd22: pixel_row = 32'b00000000011111000000000000000000;
        5'd23: pixel_row = 32'b00000000011111000000000000000000;
        5'd24: pixel_row = 32'b00000000111110000000000000000000;
        5'd25: pixel_row = 32'b00000001111100000000000000000000;
        5'd26: pixel_row = 32'b00000011111100000000000000000000;
        5'd27: pixel_row = 32'b00000011111000000000000000000000;
        5'd28: pixel_row = 32'b00000111110000000000000000000000;
        5'd29: pixel_row = 32'b00001111100000000000000000000000;
        5'd30: pixel_row = 32'b00001111000000000000000000000000;
        5'd31: pixel_row = 32'b00001100000000000000000000000000;
    endcase
end

           4'h8: begin // 8 karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00000000000011111111111100000000;
        5'd1:  pixel_row = 32'b00000000011111111111111111000000;
        5'd2:  pixel_row = 32'b00000001111111111111111111100000;
        5'd3:  pixel_row = 32'b00000011111000000000000111110000;
        5'd4:  pixel_row = 32'b00000111100000000000000011110000;
        5'd5:  pixel_row = 32'b00001111000000000000000001111000;
        5'd6:  pixel_row = 32'b00001111000000000000000001111000;
        5'd7:  pixel_row = 32'b00001110000000000000000001111000;
        5'd8:  pixel_row = 32'b00001110000000000000000001111000;
        5'd9:  pixel_row = 32'b00001111000000000000000001111000;
        5'd10: pixel_row = 32'b00001111000000000000000001111000;
        5'd11: pixel_row = 32'b00001111000000000000000011110000;
        5'd12: pixel_row = 32'b00000111100000000000000011110000;
        5'd13: pixel_row = 32'b00000011111000000000001111100000;
        5'd14: pixel_row = 32'b00000001111111111111111111000000;
        5'd15: pixel_row = 32'b00000000111111111111111110000000;
        5'd16: pixel_row = 32'b00000001111111111111111111000000;
        5'd17: pixel_row = 32'b00000011110000000000000111110000;
        5'd18: pixel_row = 32'b00000111100000000000000011111000;
        5'd19: pixel_row = 32'b00001111000000000000000001111000;
        5'd20: pixel_row = 32'b00001110000000000000000001111100;
        5'd21: pixel_row = 32'b00001110000000000000000001111100;
        5'd22: pixel_row = 32'b00001110000000000000000001111100;
        5'd23: pixel_row = 32'b00001111000000000000000001111100;
        5'd24: pixel_row = 32'b00001111000000000000000011111000;
        5'd25: pixel_row = 32'b00001111100000000000000011111000;
        5'd26: pixel_row = 32'b00000111111000000000001111110000;
        5'd27: pixel_row = 32'b00000011111111111111111111100000;
        5'd28: pixel_row = 32'b00000001111111111111111111000000;
        5'd29: pixel_row = 32'b00000000011111111111111110000000;
        5'd30: pixel_row = 32'b00000000001111111111111100000000;
        5'd31: pixel_row = 32'b00000000000001111111111000000000;
    endcase
end

            4'h9: begin // 9 karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00000000000001111111111100000000;
        5'd1:  pixel_row = 32'b00000000001111111111111111000000;
        5'd2:  pixel_row = 32'b00000000011111111111111111100000;
        5'd3:  pixel_row = 32'b00000000111110000000000111110000;
        5'd4:  pixel_row = 32'b00000001111100000000000011111000;
        5'd5:  pixel_row = 32'b00000001111000000000000001111000;
        5'd6:  pixel_row = 32'b00000011110000000000000001111000;
        5'd7:  pixel_row = 32'b00000011110000000000000001111100;
        5'd8:  pixel_row = 32'b00000111100000000000000001111100;
        5'd9:  pixel_row = 32'b00000111100000000000000001111100;
        5'd10: pixel_row = 32'b00000111100000000000000001111100;
        5'd11: pixel_row = 32'b00000111100000000000000011111100;
        5'd12: pixel_row = 32'b00000111100000000000000111111100;
        5'd13: pixel_row = 32'b00000011110000000000011111111000;
        5'd14: pixel_row = 32'b00000011111111111111111111111000;
        5'd15: pixel_row = 32'b00000001111111111111111111110000;
        5'd16: pixel_row = 32'b00000000111111111111111111110000;
        5'd17: pixel_row = 32'b00000000000000000000000011111000;
        5'd18: pixel_row = 32'b00000000000000000000000011111000;
        5'd19: pixel_row = 32'b00000000000000000000000011111000;
        5'd20: pixel_row = 32'b00000000000000000000000011111000;
        5'd21: pixel_row = 32'b00000000000000000000000011111000;
        5'd22: pixel_row = 32'b00000000000000000000000111110000;
        5'd23: pixel_row = 32'b00000000000000000000001111110000;
        5'd24: pixel_row = 32'b00000000000000000000001111110000;
        5'd25: pixel_row = 32'b00000000000000000000011111100000;
        5'd26: pixel_row = 32'b00000000000000000000011111100000;
        5'd27: pixel_row = 32'b00000000000000000000111111000000;
        5'd28: pixel_row = 32'b00000000000000000001111110000000;
        5'd29: pixel_row = 32'b00000000000000000001111100000000;
        5'd30: pixel_row = 32'b00000000000000000011111000000000;
        5'd31: pixel_row = 32'b00000000000000000011110000000000;
    endcase
end
            
           
           4'hF: begin // Bo?luk karakteri için
    case (row)
        5'd0:  pixel_row = 32'b00000000000000000000000000000000;
        5'd1:  pixel_row = 32'b00000000000000000000000000000000;
        5'd2:  pixel_row = 32'b00000000000000000000000000000000;
        5'd3:  pixel_row = 32'b00000000000000000000000000000000;
        5'd4:  pixel_row = 32'b00000000000000000000000000000000;
        5'd5:  pixel_row = 32'b00000000000000000000000000000000;
        5'd6:  pixel_row = 32'b00000000000000000000000000000000;
        5'd7:  pixel_row = 32'b00000000000000000000000000000000;
        5'd8:  pixel_row = 32'b00000000000000000000000000000000;
        5'd9:  pixel_row = 32'b00000000000000000000000000000000;
        5'd10: pixel_row = 32'b00000000000000000000000000000000;
        5'd11: pixel_row = 32'b00000000000000000000000000000000;
        5'd12: pixel_row = 32'b00000000000000000000000000000000;
        5'd13: pixel_row = 32'b00000000000000000000000000000000;
        5'd14: pixel_row = 32'b00000000000000000000000000000000;
        5'd15: pixel_row = 32'b00000000000000000000000000000000;
        5'd16: pixel_row = 32'b00000000000000000000000000000000;
        5'd17: pixel_row = 32'b00000000000000000000000000000000;
        5'd18: pixel_row = 32'b00000000000000000000000000000000;
        5'd19: pixel_row = 32'b00000000000000000000000000000000;
        5'd20: pixel_row = 32'b00000000000000000000000000000000;
        5'd21: pixel_row = 32'b00000000000000000000000000000000;
        5'd22: pixel_row = 32'b00000000000000000000000000000000;
        5'd23: pixel_row = 32'b00000000000000000000000000000000;
        5'd24: pixel_row = 32'b00000000000000000000000000000000;
        5'd25: pixel_row = 32'b00000000000000000000000000000000;
        5'd26: pixel_row = 32'b00000000000000000000000000000000;
        5'd27: pixel_row = 32'b00000000000000000000000000000000;
        5'd28: pixel_row = 32'b00000000000000000000000000000000;
        5'd29: pixel_row = 32'b00000000000000000000000000000000;
        5'd30: pixel_row = 32'b00000000000000000000000000000000;
        5'd31: pixel_row = 32'b00000000000000000000000000000000;
    endcase
end
            default: begin
                pixel_row = 8'b00000000; // Geçersiz karakter için bo? sat?r
            end
        endcase
    end
endmodule